XSpice Test

.model myclk clk (freq=10)

.model dac1 dac_bridge (out_low = 0.0
+                       out_high = 3.3
+                       out_undef = 1.7
+                       input_load = 5.0e-12
+                       t_ris e = 50e-9
+                       t_fall = 20e-9)

aclk dout myclk

abridge1 [dout] [aout] dac1

R aout 0 1k

.tran 10ms 1s

.control
pre_codemodel ./codemodel/clk.cm
run
plot v(aout) v(dout)
.endc

.end
